

-- Addition of two 5x5 matrices




-- the matrix creation is redundant (puts 1 in R0 everytime we want to put 1 into memory)
-- Just put there if we want to set different values for the matrix, if now, we should remove all x"3001" operations after the first one


--matrix 0 (columns created from left to right)(items in colums are created top to bottom)

--column 0 

0 => x"3001",			-- No. 1 -> R0
1 => x"1000",			-- R0    -> Mem[0]

2 => x"3001",			-- No. 1 -> R0
3 => x"1001",			-- R0    -> Mem[1]

4 => x"3001",			-- No. 1 -> R0
5 => x"1002",			-- R0    -> Mem[2]

6 => x"3001",			-- No. 1 -> R0
7 => x"1003",			-- R0    -> Mem[3]

8 => x"3001",			-- No. 1 -> R0
9 => x"1004",			-- R0    -> Mem[4]

--column 1

10 => x"3001",			-- No. 1 -> R0
11 => x"1005",			-- R0    -> Mem[5]

12 => x"3001",			-- No. 1 -> R0
13 => x"1006",			-- R0    -> Mem[6]

14 => x"3001",			-- No. 1 -> R0
15 => x"1007",			-- R0    -> Mem[7]

16 => x"3001",			-- No. 1 -> R0
17 => x"1008",			-- R0    -> Mem[8]

18 => x"3001",			-- No. 1 -> R0
19 => x"1009",			-- R0    -> Mem[9]

--column 2

20 => x"3001",			-- No. 1 -> R0
21 => x"100A",			-- R0    -> Mem[10]

22 => x"3001",			-- No. 1 -> R0
23 => x"100B",			-- R0    -> Mem[11]

24 => x"3001",			-- No. 1 -> R0
25 => x"100C",			-- R0    -> Mem[12]

26 => x"3001",			-- No. 1 -> R0
27 => x"100D",			-- R0    -> Mem[13]

28 => x"3001",			-- No. 1 -> R0
29 => x"100E",			-- R0    -> Mem[14]

--column 3

30 => x"3001",			-- No. 1 -> R0
31 => x"100F",			-- R0    -> Mem[15]

32 => x"3001",			-- No. 1 -> R0
33 => x"1010",			-- R0    -> Mem[16]

34 => x"3001",			-- No. 1 -> R0
35 => x"1011",			-- R0    -> Mem[17]

36 => x"3001",			-- No. 1 -> R0
37 => x"1012",			-- R0    -> Mem[18]

38 => x"3001",			-- No. 1 -> R0
39 => x"1013",			-- R0    -> Mem[19]

--column 4

40 => x"3001",			-- No. 1 -> R0
41 => x"1014",			-- R0    -> Mem[20]

42 => x"3001",			-- No. 1 -> R0
43 => x"1015",			-- R0    -> Mem[21]

44 => x"3001",			-- No. 1 -> R0
45 => x"1016",			-- R0    -> Mem[22]

46 => x"3001",			-- No. 1 -> R0
47 => x"1017",			-- R0    -> Mem[23]

48 => x"3001",			-- No. 1 -> R0
49 => x"1018",			-- R0    -> Mem[24]



--matrix 1


--column 0

50 => x"3001",			-- No. 1 -> R0
51 => x"1019",			-- R0    -> Mem[25]

52 => x"3001",			-- No. 1 -> R0
53 => x"101A",			-- R0    -> Mem[26]

54 => x"3001",			-- No. 1 -> R0
55 => x"101B",			-- R0    -> Mem[27]

56 => x"3001",			-- No. 1 -> R0
57 => x"101C",			-- R0    -> Mem[28]

58 => x"3001",			-- No. 1 -> R0
59 => x"101D",			-- R0    -> Mem[29]

--column 1

60 => x"3001",			-- No. 1 -> R0
61 => x"101E",			-- R0    -> Mem[30]

62 => x"3001",			-- No. 1 -> R0
63 => x"101F",			-- R0    -> Mem[31]

64 => x"3001",			-- No. 1 -> R0
65 => x"1020",			-- R0    -> Mem[32]

66 => x"3001",			-- No. 1 -> R0
67 => x"1021",			-- R0    -> Mem[33]

68 => x"3001",			-- No. 1 -> R0
69 => x"1022",			-- R0    -> Mem[34]

--column 2

70 => x"3001",			-- No. 1 -> R0
71 => x"1023",			-- R0    -> Mem[35]

72 => x"3001",			-- No. 1 -> R0
73 => x"1024",			-- R0    -> Mem[36]

74 => x"3001",			-- No. 1 -> R0
75 => x"1025",			-- R0    -> Mem[37]

76 => x"3001",			-- No. 1 -> R0
77 => x"1026",			-- R0    -> Mem[38]

78 => x"3001",			-- No. 1 -> R0
79 => x"1027",			-- R0    -> Mem[39]

--column 3

80 => x"3001",			-- No. 1 -> R0
81 => x"1028",			-- R0    -> Mem[40]

82 => x"3001",			-- No. 1 -> R0
83 => x"1029",			-- R0    -> Mem[41]

84 => x"3001",			-- No. 1 -> R0
85 => x"102A",			-- R0    -> Mem[42]

86 => x"3001",			-- No. 1 -> R0
87 => x"102B",			-- R0    -> Mem[43]

88 => x"3001",			-- No. 1 -> R0
89 => x"102C",			-- R0    -> Mem[44]

--column 4

90 => x"3001",			-- No. 1 -> R0
91 => x"102D",			-- R0    -> Mem[45]

92 => x"3001",			-- No. 1 -> R0
93 => x"102E",			-- R0    -> Mem[46]

94 => x"3001",			-- No. 1 -> R0
95 => x"102F",			-- R0    -> Mem[47]

96 => x"3001",			-- No. 1 -> R0
97 => x"1030",			-- R0    -> Mem[48]

98 => x"3001",			-- No. 1 -> R0
99 => x"1031",			-- R0    -> Mem[49]






-- matrix addition. result found in memory location mem[50]..mem[74]
		(starts adding from top left corner then goes top-down following the columns)


100 => x"0000",			-- Mem[0] -> R0
101 => x"0119",			-- Mem[25]-> R1
102 => x"4010",			-- R0 	   = R0 + R1
103 => x"1032",			-- R0     -> Mem[50]

104 => x"0001",			-- Mem[1] -> R0
105 => x"011A",			-- Mem[26]-> R1
106 => x"4010",			-- R0 	   = R0 + R1
107 => x"1033",			-- R0     -> Mem[51]

108 => x"0002",			-- Mem[2] -> R0
109 => x"011B",			-- Mem[27]-> R1
110 => x"4010",			-- R0 	   = R0 + R1
111 => x"1034",			-- R0     -> Mem[52]

112 => x"0003",			-- Mem[3] -> R0
113 => x"011C",			-- Mem[28]-> R1
114 => x"4010",			-- R0 	   = R0 + R1
115 => x"1035",			-- R0     -> Mem[53]

116 => x"0004",			-- Mem[4] -> R0
117 => x"011D",			-- Mem[29]-> R1
118 => x"4010",			-- R0 	   = R0 + R1
119 => x"1036",			-- R0     -> Mem[54]




120 => x"0005",			-- Mem[5] -> R0
121 => x"011E",			-- Mem[30]-> R1
122 => x"4010",			-- R0 	   = R0 + R1
123 => x"1037",			-- R0     -> Mem[55]

124 => x"0006",			-- Mem[6] -> R0
125 => x"011F",			-- Mem[31]-> R1
126 => x"4010",			-- R0 	   = R0 + R1
127 => x"1038",			-- R0     -> Mem[56]

128 => x"0007",			-- Mem[7] -> R0
129 => x"0120",			-- Mem[32]-> R1
130 => x"4010",			-- R0 	   = R0 + R1
131 => x"1039",			-- R0     -> Mem[57]

132 => x"0008",			-- Mem[8] -> R0
133 => x"0121",			-- Mem[33]-> R1
134 => x"4010",			-- R0 	   = R0 + R1
135 => x"103A",			-- R0     -> Mem[58]

136 => x"0009",			-- Mem[9] -> R0
137 => x"0122",			-- Mem[34]-> R1
138 => x"4010",			-- R0 	   = R0 + R1
139 => x"103B",			-- R0     -> Mem[59]




140 => x"000A",			-- Mem[10]-> R0
141 => x"0123",			-- Mem[35]-> R1
142 => x"4010",			-- R0 	   = R0 + R1
143 => x"103C",			-- R0     -> Mem[60]

144 => x"000B",			-- Mem[11] -> R0
145 => x"0124",			-- Mem[36]-> R1
146 => x"4010",			-- R0 	   = R0 + R1
147 => x"103D",			-- R0     -> Mem[61]

148 => x"000C",			-- Mem[12] -> R0
149 => x"0125",			-- Mem[37]-> R1
150 => x"4010",			-- R0 	   = R0 + R1
151 => x"103E",			-- R0     -> Mem[62]

152 => x"000D",			-- Mem[13] -> R0
153 => x"0126",			-- Mem[38]-> R1
154 => x"4010",			-- R0 	   = R0 + R1
155 => x"103F",			-- R0     -> Mem[63]

156 => x"000E",			-- Mem[14] -> R0
157 => x"0127",			-- Mem[39]-> R1
158 => x"4010",			-- R0 	   = R0 + R1
159 => x"1040", 		-- R0     -> Mem[64]




160 => x"000F",			-- Mem[15] -> R0
161 => x"0128",			-- Mem[40]-> R1
162 => x"4010",			-- R0 	   = R0 + R1
163 => x"1041",			-- R0     -> Mem[65]

164 => x"0010",			-- Mem[16] -> R0
165 => x"0129",			-- Mem[41]-> R1
166 => x"4010",			-- R0 	   = R0 + R1
167 => x"1042",			-- R0     -> Mem[66]

168 => x"0011",			-- Mem[17] -> R0
169 => x"012A",			-- Mem[42]-> R1
170 => x"4010",			-- R0 	   = R0 + R1
171 => x"1043",			-- R0     -> Mem[67]

172 => x"0012",			-- Mem[18] -> R0
173 => x"012B",			-- Mem[43]-> R1
174 => x"4010",			-- R0 	   = R0 + R1
175 => x"1044",			-- R0     -> Mem[68]

176 => x"0013",			-- Mem[19] -> R0
177 => x"012C",			-- Mem[44]-> R1
178 => x"4010",			-- R0 	   = R0 + R1
179 => x"1045",			-- R0     -> Mem[69]




180 => x"0014",			-- Mem[20] -> R0
181 => x"012D",			-- Mem[45]-> R1
182 => x"4010",			-- R0 	   = R0 + R1
183 => x"1046",			-- R0     -> Mem[70]

184 => x"0015",			-- Mem[21] -> R0
185 => x"012E",			-- Mem[46]-> R1
186 => x"4010",			-- R0 	   = R0 + R1
187 => x"1047",			-- R0     -> Mem[71]

188 => x"0016",			-- Mem[22] -> R0
189 => x"012F",			-- Mem[47]-> R1
190 => x"4010",			-- R0 	   = R0 + R1
191 => x"1048",			-- R0     -> Mem[72]

192 => x"0017",			-- Mem[23] -> R0
193 => x"0130",			-- Mem[48]-> R1
194 => x"4010",			-- R0 	   = R0 + R1
195 => x"1049",			-- R0     -> Mem[73]

196 => x"0018",			-- Mem[24] -> R0
197 => x"0131",			-- Mem[49]-> R1
198 => x"4010",			-- R0 	   = R0 + R1
199 => x"104A",			-- R0     -> Mem[74]






