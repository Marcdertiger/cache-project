
--------------------------------------------------------
-- Simple Microprocessor Design 
--
-- alu has functions of bypass, addition and subtraction
-- alu.vhd
--------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;  
use work.MP_lib.all;

-- addition of logic to compare if a register is of value 25 decimal.
-- allows for 5x5 matrix operations.

-- future implementation may include comparism to any number, more complex
-- logic is needed to do so. Not necessary for the limited use of such logic.


entity alu is
port (	num_A: 	in std_logic_vector(15 downto 0);
		num_B: 	in std_logic_vector(15 downto 0);
		jpsign:	in std_logic;						 -- JMP?	
		ALUs:	in std_logic_vector(1 downto 0);     -- OP selector
		ALUz:	out std_logic;                       -- Reached 0!   
		ALUout:	out std_logic_vector(15 downto 0);    -- final calc value
		jpsign2:	in std_logic						 -- JMP2
);
end alu;

architecture behv of alu is

signal alu_tmp: std_logic_vector(15 downto 0);

begin

	process(num_A, num_B, ALUs)
	begin			
		case ALUs is
		  when "00" => alu_tmp <= num_A;
		  when "01" => alu_tmp <= num_B;
		  when "10" => alu_tmp <= num_A + num_B;
		  when "11" => alu_tmp <= num_A - num_B;
		  when others =>
	    end case; 					  
	end process;
	
	process(jpsign, alu_tmp,jpsign2)
	begin
	
	--for some reason, jz2 jumps all the time
		if (jpsign = '1' and alu_tmp = ZERO)or(jpsign2 = '1' and (alu_tmp > ZERO)) then
			ALUz <= '1';
		else
			ALUz <= '0';
		end if;
		
		--if (jpsign2 = '1' and alu_tmp /= ZERO) then
		--	ALUz <= '1';
		--else
		--	ALUz <= '0';
		--end if;
	end process;					
	
	ALUout <= alu_tmp;
	
end behv;









