-- SRAM

-- contains the data lines of the cache

-- 8 lined of 4 words, words of 16 bits